package ahb2apb_pkg;

//`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "uvm_macros.svh"

//included files of all the components that I have created
`include "ahb2apb_transaction.sv"
`include "ahb2apb_base_seq.sv"
`include "ahb2apb_write_seq.sv"
`include "ahb2apb_single_seq.sv"
`include "ahb2apb_incr_seq.sv"
`include "ahb2apb_incr4_seq.sv"
`include "ahb2apb_incr8_seq.sv"
`include "ahb2apb_incr16_seq.sv"
`include "ahb2apb_wrap4_seq.sv"
`include "ahb2apb_wrap8_seq.sv"
`include "ahb2apb_wrap16_seq.sv"
`include "ahb2apb_master_sequencer.sv"
`include "ahb2apb_master_driver.sv"
`include "ahb2apb_slave_driver.sv"
`include "ahb2apb_master_monitor.sv"
`include "ahb2apb_slave_monitor.sv"
`include "ahb2apb_master_agent.sv"
`include "ahb2apb_slave_agent.sv"
`include "ahb2apb_scoreboard.sv"
`include "ahb2apb_subscriber.sv"
`include "ahb2apb_env.sv"
`include "ahb2apb_base_test.sv"
`include "ahb2apb_test.sv"
`include "ahb2apb_single_test.sv"
`include "ahb2apb_incr_test.sv"
`include "ahb2apb_wrap_test.sv"


endpackage
